module rom(input [4:0] n1, input [4:0] n2, output [9:0] res);

    reg [9:0] rom [1023:0];

    initial
    begin

        rom[0] = 10'b0000000000; // 0 * 0 = 0
        rom[1] = 10'b0000000000; // 0 * 1 = 0
        rom[2] = 10'b0000000000; // 0 * 2 = 0
        rom[3] = 10'b0000000000; // 0 * 3 = 0
        rom[4] = 10'b0000000000; // 0 * 4 = 0
        rom[5] = 10'b0000000000; // 0 * 5 = 0
        rom[6] = 10'b0000000000; // 0 * 6 = 0
        rom[7] = 10'b0000000000; // 0 * 7 = 0
        rom[8] = 10'b0000000000; // 0 * 8 = 0
        rom[9] = 10'b0000000000; // 0 * 9 = 0
        rom[10] = 10'b0000000000; // 0 * 10 = 0
        rom[11] = 10'b0000000000; // 0 * 11 = 0
        rom[12] = 10'b0000000000; // 0 * 12 = 0
        rom[13] = 10'b0000000000; // 0 * 13 = 0
        rom[14] = 10'b0000000000; // 0 * 14 = 0
        rom[15] = 10'b0000000000; // 0 * 15 = 0
        rom[16] = 10'b0000000000; // 0 * 16 = 0
        rom[17] = 10'b0000000000; // 0 * 17 = 0
        rom[18] = 10'b0000000000; // 0 * 18 = 0
        rom[19] = 10'b0000000000; // 0 * 19 = 0
        rom[20] = 10'b0000000000; // 0 * 20 = 0
        rom[21] = 10'b0000000000; // 0 * 21 = 0
        rom[22] = 10'b0000000000; // 0 * 22 = 0
        rom[23] = 10'b0000000000; // 0 * 23 = 0
        rom[24] = 10'b0000000000; // 0 * 24 = 0
        rom[25] = 10'b0000000000; // 0 * 25 = 0
        rom[26] = 10'b0000000000; // 0 * 26 = 0
        rom[27] = 10'b0000000000; // 0 * 27 = 0
        rom[28] = 10'b0000000000; // 0 * 28 = 0
        rom[29] = 10'b0000000000; // 0 * 29 = 0
        rom[30] = 10'b0000000000; // 0 * 30 = 0
        rom[31] = 10'b0000000000; // 0 * 31 = 0
        rom[32] = 10'b0000000000; // 1 * 0 = 0
        rom[33] = 10'b0000000001; // 1 * 1 = 1
        rom[34] = 10'b0000000010; // 1 * 2 = 2
        rom[35] = 10'b0000000011; // 1 * 3 = 3
        rom[36] = 10'b0000000100; // 1 * 4 = 4
        rom[37] = 10'b0000000101; // 1 * 5 = 5
        rom[38] = 10'b0000000110; // 1 * 6 = 6
        rom[39] = 10'b0000000111; // 1 * 7 = 7
        rom[40] = 10'b0000001000; // 1 * 8 = 8
        rom[41] = 10'b0000001001; // 1 * 9 = 9
        rom[42] = 10'b0000001010; // 1 * 10 = 10
        rom[43] = 10'b0000001011; // 1 * 11 = 11
        rom[44] = 10'b0000001100; // 1 * 12 = 12
        rom[45] = 10'b0000001101; // 1 * 13 = 13
        rom[46] = 10'b0000001110; // 1 * 14 = 14
        rom[47] = 10'b0000001111; // 1 * 15 = 15
        rom[48] = 10'b0000010000; // 1 * 16 = 16
        rom[49] = 10'b0000010001; // 1 * 17 = 17
        rom[50] = 10'b0000010010; // 1 * 18 = 18
        rom[51] = 10'b0000010011; // 1 * 19 = 19
        rom[52] = 10'b0000010100; // 1 * 20 = 20
        rom[53] = 10'b0000010101; // 1 * 21 = 21
        rom[54] = 10'b0000010110; // 1 * 22 = 22
        rom[55] = 10'b0000010111; // 1 * 23 = 23
        rom[56] = 10'b0000011000; // 1 * 24 = 24
        rom[57] = 10'b0000011001; // 1 * 25 = 25
        rom[58] = 10'b0000011010; // 1 * 26 = 26
        rom[59] = 10'b0000011011; // 1 * 27 = 27
        rom[60] = 10'b0000011100; // 1 * 28 = 28
        rom[61] = 10'b0000011101; // 1 * 29 = 29
        rom[62] = 10'b0000011110; // 1 * 30 = 30
        rom[63] = 10'b0000011111; // 1 * 31 = 31
        rom[64] = 10'b0000000000; // 2 * 0 = 0
        rom[65] = 10'b0000000010; // 2 * 1 = 2
        rom[66] = 10'b0000000100; // 2 * 2 = 4
        rom[67] = 10'b0000000110; // 2 * 3 = 6
        rom[68] = 10'b0000001000; // 2 * 4 = 8
        rom[69] = 10'b0000001010; // 2 * 5 = 10
        rom[70] = 10'b0000001100; // 2 * 6 = 12
        rom[71] = 10'b0000001110; // 2 * 7 = 14
        rom[72] = 10'b0000010000; // 2 * 8 = 16
        rom[73] = 10'b0000010010; // 2 * 9 = 18
        rom[74] = 10'b0000010100; // 2 * 10 = 20
        rom[75] = 10'b0000010110; // 2 * 11 = 22
        rom[76] = 10'b0000011000; // 2 * 12 = 24
        rom[77] = 10'b0000011010; // 2 * 13 = 26
        rom[78] = 10'b0000011100; // 2 * 14 = 28
        rom[79] = 10'b0000011110; // 2 * 15 = 30
        rom[80] = 10'b0000100000; // 2 * 16 = 32
        rom[81] = 10'b0000100010; // 2 * 17 = 34
        rom[82] = 10'b0000100100; // 2 * 18 = 36
        rom[83] = 10'b0000100110; // 2 * 19 = 38
        rom[84] = 10'b0000101000; // 2 * 20 = 40
        rom[85] = 10'b0000101010; // 2 * 21 = 42
        rom[86] = 10'b0000101100; // 2 * 22 = 44
        rom[87] = 10'b0000101110; // 2 * 23 = 46
        rom[88] = 10'b0000110000; // 2 * 24 = 48
        rom[89] = 10'b0000110010; // 2 * 25 = 50
        rom[90] = 10'b0000110100; // 2 * 26 = 52
        rom[91] = 10'b0000110110; // 2 * 27 = 54
        rom[92] = 10'b0000111000; // 2 * 28 = 56
        rom[93] = 10'b0000111010; // 2 * 29 = 58
        rom[94] = 10'b0000111100; // 2 * 30 = 60
        rom[95] = 10'b0000111110; // 2 * 31 = 62
        rom[96] = 10'b0000000000; // 3 * 0 = 0
        rom[97] = 10'b0000000011; // 3 * 1 = 3
        rom[98] = 10'b0000000110; // 3 * 2 = 6
        rom[99] = 10'b0000001001; // 3 * 3 = 9
        rom[100] = 10'b0000001100; // 3 * 4 = 12
        rom[101] = 10'b0000001111; // 3 * 5 = 15
        rom[102] = 10'b0000010010; // 3 * 6 = 18
        rom[103] = 10'b0000010101; // 3 * 7 = 21
        rom[104] = 10'b0000011000; // 3 * 8 = 24
        rom[105] = 10'b0000011011; // 3 * 9 = 27
        rom[106] = 10'b0000011110; // 3 * 10 = 30
        rom[107] = 10'b0000100001; // 3 * 11 = 33
        rom[108] = 10'b0000100100; // 3 * 12 = 36
        rom[109] = 10'b0000100111; // 3 * 13 = 39
        rom[110] = 10'b0000101010; // 3 * 14 = 42
        rom[111] = 10'b0000101101; // 3 * 15 = 45
        rom[112] = 10'b0000110000; // 3 * 16 = 48
        rom[113] = 10'b0000110011; // 3 * 17 = 51
        rom[114] = 10'b0000110110; // 3 * 18 = 54
        rom[115] = 10'b0000111001; // 3 * 19 = 57
        rom[116] = 10'b0000111100; // 3 * 20 = 60
        rom[117] = 10'b0000111111; // 3 * 21 = 63
        rom[118] = 10'b0001000010; // 3 * 22 = 66
        rom[119] = 10'b0001000101; // 3 * 23 = 69
        rom[120] = 10'b0001001000; // 3 * 24 = 72
        rom[121] = 10'b0001001011; // 3 * 25 = 75
        rom[122] = 10'b0001001110; // 3 * 26 = 78
        rom[123] = 10'b0001010001; // 3 * 27 = 81
        rom[124] = 10'b0001010100; // 3 * 28 = 84
        rom[125] = 10'b0001010111; // 3 * 29 = 87
        rom[126] = 10'b0001011010; // 3 * 30 = 90
        rom[127] = 10'b0001011101; // 3 * 31 = 93
        rom[128] = 10'b0000000000; // 4 * 0 = 0
        rom[129] = 10'b0000000100; // 4 * 1 = 4
        rom[130] = 10'b0000001000; // 4 * 2 = 8
        rom[131] = 10'b0000001100; // 4 * 3 = 12
        rom[132] = 10'b0000010000; // 4 * 4 = 16
        rom[133] = 10'b0000010100; // 4 * 5 = 20
        rom[134] = 10'b0000011000; // 4 * 6 = 24
        rom[135] = 10'b0000011100; // 4 * 7 = 28
        rom[136] = 10'b0000100000; // 4 * 8 = 32
        rom[137] = 10'b0000100100; // 4 * 9 = 36
        rom[138] = 10'b0000101000; // 4 * 10 = 40
        rom[139] = 10'b0000101100; // 4 * 11 = 44
        rom[140] = 10'b0000110000; // 4 * 12 = 48
        rom[141] = 10'b0000110100; // 4 * 13 = 52
        rom[142] = 10'b0000111000; // 4 * 14 = 56
        rom[143] = 10'b0000111100; // 4 * 15 = 60
        rom[144] = 10'b0001000000; // 4 * 16 = 64
        rom[145] = 10'b0001000100; // 4 * 17 = 68
        rom[146] = 10'b0001001000; // 4 * 18 = 72
        rom[147] = 10'b0001001100; // 4 * 19 = 76
        rom[148] = 10'b0001010000; // 4 * 20 = 80
        rom[149] = 10'b0001010100; // 4 * 21 = 84
        rom[150] = 10'b0001011000; // 4 * 22 = 88
        rom[151] = 10'b0001011100; // 4 * 23 = 92
        rom[152] = 10'b0001100000; // 4 * 24 = 96
        rom[153] = 10'b0001100100; // 4 * 25 = 100
        rom[154] = 10'b0001101000; // 4 * 26 = 104
        rom[155] = 10'b0001101100; // 4 * 27 = 108
        rom[156] = 10'b0001110000; // 4 * 28 = 112
        rom[157] = 10'b0001110100; // 4 * 29 = 116
        rom[158] = 10'b0001111000; // 4 * 30 = 120
        rom[159] = 10'b0001111100; // 4 * 31 = 124
        rom[160] = 10'b0000000000; // 5 * 0 = 0
        rom[161] = 10'b0000000101; // 5 * 1 = 5
        rom[162] = 10'b0000001010; // 5 * 2 = 10
        rom[163] = 10'b0000001111; // 5 * 3 = 15
        rom[164] = 10'b0000010100; // 5 * 4 = 20
        rom[165] = 10'b0000011001; // 5 * 5 = 25
        rom[166] = 10'b0000011110; // 5 * 6 = 30
        rom[167] = 10'b0000100011; // 5 * 7 = 35
        rom[168] = 10'b0000101000; // 5 * 8 = 40
        rom[169] = 10'b0000101101; // 5 * 9 = 45
        rom[170] = 10'b0000110010; // 5 * 10 = 50
        rom[171] = 10'b0000110111; // 5 * 11 = 55
        rom[172] = 10'b0000111100; // 5 * 12 = 60
        rom[173] = 10'b0001000001; // 5 * 13 = 65
        rom[174] = 10'b0001000110; // 5 * 14 = 70
        rom[175] = 10'b0001001011; // 5 * 15 = 75
        rom[176] = 10'b0001010000; // 5 * 16 = 80
        rom[177] = 10'b0001010101; // 5 * 17 = 85
        rom[178] = 10'b0001011010; // 5 * 18 = 90
        rom[179] = 10'b0001011111; // 5 * 19 = 95
        rom[180] = 10'b0001100100; // 5 * 20 = 100
        rom[181] = 10'b0001101001; // 5 * 21 = 105
        rom[182] = 10'b0001101110; // 5 * 22 = 110
        rom[183] = 10'b0001110011; // 5 * 23 = 115
        rom[184] = 10'b0001111000; // 5 * 24 = 120
        rom[185] = 10'b0001111101; // 5 * 25 = 125
        rom[186] = 10'b0010000010; // 5 * 26 = 130
        rom[187] = 10'b0010000111; // 5 * 27 = 135
        rom[188] = 10'b0010001100; // 5 * 28 = 140
        rom[189] = 10'b0010010001; // 5 * 29 = 145
        rom[190] = 10'b0010010110; // 5 * 30 = 150
        rom[191] = 10'b0010011011; // 5 * 31 = 155
        rom[192] = 10'b0000000000; // 6 * 0 = 0
        rom[193] = 10'b0000000110; // 6 * 1 = 6
        rom[194] = 10'b0000001100; // 6 * 2 = 12
        rom[195] = 10'b0000010010; // 6 * 3 = 18
        rom[196] = 10'b0000011000; // 6 * 4 = 24
        rom[197] = 10'b0000011110; // 6 * 5 = 30
        rom[198] = 10'b0000100100; // 6 * 6 = 36
        rom[199] = 10'b0000101010; // 6 * 7 = 42
        rom[200] = 10'b0000110000; // 6 * 8 = 48
        rom[201] = 10'b0000110110; // 6 * 9 = 54
        rom[202] = 10'b0000111100; // 6 * 10 = 60
        rom[203] = 10'b0001000010; // 6 * 11 = 66
        rom[204] = 10'b0001001000; // 6 * 12 = 72
        rom[205] = 10'b0001001110; // 6 * 13 = 78
        rom[206] = 10'b0001010100; // 6 * 14 = 84
        rom[207] = 10'b0001011010; // 6 * 15 = 90
        rom[208] = 10'b0001100000; // 6 * 16 = 96
        rom[209] = 10'b0001100110; // 6 * 17 = 102
        rom[210] = 10'b0001101100; // 6 * 18 = 108
        rom[211] = 10'b0001110010; // 6 * 19 = 114
        rom[212] = 10'b0001111000; // 6 * 20 = 120
        rom[213] = 10'b0001111110; // 6 * 21 = 126
        rom[214] = 10'b0010000100; // 6 * 22 = 132
        rom[215] = 10'b0010001010; // 6 * 23 = 138
        rom[216] = 10'b0010010000; // 6 * 24 = 144
        rom[217] = 10'b0010010110; // 6 * 25 = 150
        rom[218] = 10'b0010011100; // 6 * 26 = 156
        rom[219] = 10'b0010100010; // 6 * 27 = 162
        rom[220] = 10'b0010101000; // 6 * 28 = 168
        rom[221] = 10'b0010101110; // 6 * 29 = 174
        rom[222] = 10'b0010110100; // 6 * 30 = 180
        rom[223] = 10'b0010111010; // 6 * 31 = 186
        rom[224] = 10'b0000000000; // 7 * 0 = 0
        rom[225] = 10'b0000000111; // 7 * 1 = 7
        rom[226] = 10'b0000001110; // 7 * 2 = 14
        rom[227] = 10'b0000010101; // 7 * 3 = 21
        rom[228] = 10'b0000011100; // 7 * 4 = 28
        rom[229] = 10'b0000100011; // 7 * 5 = 35
        rom[230] = 10'b0000101010; // 7 * 6 = 42
        rom[231] = 10'b0000110001; // 7 * 7 = 49
        rom[232] = 10'b0000111000; // 7 * 8 = 56
        rom[233] = 10'b0000111111; // 7 * 9 = 63
        rom[234] = 10'b0001000110; // 7 * 10 = 70
        rom[235] = 10'b0001001101; // 7 * 11 = 77
        rom[236] = 10'b0001010100; // 7 * 12 = 84
        rom[237] = 10'b0001011011; // 7 * 13 = 91
        rom[238] = 10'b0001100010; // 7 * 14 = 98
        rom[239] = 10'b0001101001; // 7 * 15 = 105
        rom[240] = 10'b0001110000; // 7 * 16 = 112
        rom[241] = 10'b0001110111; // 7 * 17 = 119
        rom[242] = 10'b0001111110; // 7 * 18 = 126
        rom[243] = 10'b0010000101; // 7 * 19 = 133
        rom[244] = 10'b0010001100; // 7 * 20 = 140
        rom[245] = 10'b0010010011; // 7 * 21 = 147
        rom[246] = 10'b0010011010; // 7 * 22 = 154
        rom[247] = 10'b0010100001; // 7 * 23 = 161
        rom[248] = 10'b0010101000; // 7 * 24 = 168
        rom[249] = 10'b0010101111; // 7 * 25 = 175
        rom[250] = 10'b0010110110; // 7 * 26 = 182
        rom[251] = 10'b0010111101; // 7 * 27 = 189
        rom[252] = 10'b0011000100; // 7 * 28 = 196
        rom[253] = 10'b0011001011; // 7 * 29 = 203
        rom[254] = 10'b0011010010; // 7 * 30 = 210
        rom[255] = 10'b0011011001; // 7 * 31 = 217
        rom[256] = 10'b0000000000; // 8 * 0 = 0
        rom[257] = 10'b0000001000; // 8 * 1 = 8
        rom[258] = 10'b0000010000; // 8 * 2 = 16
        rom[259] = 10'b0000011000; // 8 * 3 = 24
        rom[260] = 10'b0000100000; // 8 * 4 = 32
        rom[261] = 10'b0000101000; // 8 * 5 = 40
        rom[262] = 10'b0000110000; // 8 * 6 = 48
        rom[263] = 10'b0000111000; // 8 * 7 = 56
        rom[264] = 10'b0001000000; // 8 * 8 = 64
        rom[265] = 10'b0001001000; // 8 * 9 = 72
        rom[266] = 10'b0001010000; // 8 * 10 = 80
        rom[267] = 10'b0001011000; // 8 * 11 = 88
        rom[268] = 10'b0001100000; // 8 * 12 = 96
        rom[269] = 10'b0001101000; // 8 * 13 = 104
        rom[270] = 10'b0001110000; // 8 * 14 = 112
        rom[271] = 10'b0001111000; // 8 * 15 = 120
        rom[272] = 10'b0010000000; // 8 * 16 = 128
        rom[273] = 10'b0010001000; // 8 * 17 = 136
        rom[274] = 10'b0010010000; // 8 * 18 = 144
        rom[275] = 10'b0010011000; // 8 * 19 = 152
        rom[276] = 10'b0010100000; // 8 * 20 = 160
        rom[277] = 10'b0010101000; // 8 * 21 = 168
        rom[278] = 10'b0010110000; // 8 * 22 = 176
        rom[279] = 10'b0010111000; // 8 * 23 = 184
        rom[280] = 10'b0011000000; // 8 * 24 = 192
        rom[281] = 10'b0011001000; // 8 * 25 = 200
        rom[282] = 10'b0011010000; // 8 * 26 = 208
        rom[283] = 10'b0011011000; // 8 * 27 = 216
        rom[284] = 10'b0011100000; // 8 * 28 = 224
        rom[285] = 10'b0011101000; // 8 * 29 = 232
        rom[286] = 10'b0011110000; // 8 * 30 = 240
        rom[287] = 10'b0011111000; // 8 * 31 = 248
        rom[288] = 10'b0000000000; // 9 * 0 = 0
        rom[289] = 10'b0000001001; // 9 * 1 = 9
        rom[290] = 10'b0000010010; // 9 * 2 = 18
        rom[291] = 10'b0000011011; // 9 * 3 = 27
        rom[292] = 10'b0000100100; // 9 * 4 = 36
        rom[293] = 10'b0000101101; // 9 * 5 = 45
        rom[294] = 10'b0000110110; // 9 * 6 = 54
        rom[295] = 10'b0000111111; // 9 * 7 = 63
        rom[296] = 10'b0001001000; // 9 * 8 = 72
        rom[297] = 10'b0001010001; // 9 * 9 = 81
        rom[298] = 10'b0001011010; // 9 * 10 = 90
        rom[299] = 10'b0001100011; // 9 * 11 = 99
        rom[300] = 10'b0001101100; // 9 * 12 = 108
        rom[301] = 10'b0001110101; // 9 * 13 = 117
        rom[302] = 10'b0001111110; // 9 * 14 = 126
        rom[303] = 10'b0010000111; // 9 * 15 = 135
        rom[304] = 10'b0010010000; // 9 * 16 = 144
        rom[305] = 10'b0010011001; // 9 * 17 = 153
        rom[306] = 10'b0010100010; // 9 * 18 = 162
        rom[307] = 10'b0010101011; // 9 * 19 = 171
        rom[308] = 10'b0010110100; // 9 * 20 = 180
        rom[309] = 10'b0010111101; // 9 * 21 = 189
        rom[310] = 10'b0011000110; // 9 * 22 = 198
        rom[311] = 10'b0011001111; // 9 * 23 = 207
        rom[312] = 10'b0011011000; // 9 * 24 = 216
        rom[313] = 10'b0011100001; // 9 * 25 = 225
        rom[314] = 10'b0011101010; // 9 * 26 = 234
        rom[315] = 10'b0011110011; // 9 * 27 = 243
        rom[316] = 10'b0011111100; // 9 * 28 = 252
        rom[317] = 10'b0100000101; // 9 * 29 = 261
        rom[318] = 10'b0100001110; // 9 * 30 = 270
        rom[319] = 10'b0100010111; // 9 * 31 = 279
        rom[320] = 10'b0000000000; // 10 * 0 = 0
        rom[321] = 10'b0000001010; // 10 * 1 = 10
        rom[322] = 10'b0000010100; // 10 * 2 = 20
        rom[323] = 10'b0000011110; // 10 * 3 = 30
        rom[324] = 10'b0000101000; // 10 * 4 = 40
        rom[325] = 10'b0000110010; // 10 * 5 = 50
        rom[326] = 10'b0000111100; // 10 * 6 = 60
        rom[327] = 10'b0001000110; // 10 * 7 = 70
        rom[328] = 10'b0001010000; // 10 * 8 = 80
        rom[329] = 10'b0001011010; // 10 * 9 = 90
        rom[330] = 10'b0001100100; // 10 * 10 = 100
        rom[331] = 10'b0001101110; // 10 * 11 = 110
        rom[332] = 10'b0001111000; // 10 * 12 = 120
        rom[333] = 10'b0010000010; // 10 * 13 = 130
        rom[334] = 10'b0010001100; // 10 * 14 = 140
        rom[335] = 10'b0010010110; // 10 * 15 = 150
        rom[336] = 10'b0010100000; // 10 * 16 = 160
        rom[337] = 10'b0010101010; // 10 * 17 = 170
        rom[338] = 10'b0010110100; // 10 * 18 = 180
        rom[339] = 10'b0010111110; // 10 * 19 = 190
        rom[340] = 10'b0011001000; // 10 * 20 = 200
        rom[341] = 10'b0011010010; // 10 * 21 = 210
        rom[342] = 10'b0011011100; // 10 * 22 = 220
        rom[343] = 10'b0011100110; // 10 * 23 = 230
        rom[344] = 10'b0011110000; // 10 * 24 = 240
        rom[345] = 10'b0011111010; // 10 * 25 = 250
        rom[346] = 10'b0100000100; // 10 * 26 = 260
        rom[347] = 10'b0100001110; // 10 * 27 = 270
        rom[348] = 10'b0100011000; // 10 * 28 = 280
        rom[349] = 10'b0100100010; // 10 * 29 = 290
        rom[350] = 10'b0100101100; // 10 * 30 = 300
        rom[351] = 10'b0100110110; // 10 * 31 = 310
        rom[352] = 10'b0000000000; // 11 * 0 = 0
        rom[353] = 10'b0000001011; // 11 * 1 = 11
        rom[354] = 10'b0000010110; // 11 * 2 = 22
        rom[355] = 10'b0000100001; // 11 * 3 = 33
        rom[356] = 10'b0000101100; // 11 * 4 = 44
        rom[357] = 10'b0000110111; // 11 * 5 = 55
        rom[358] = 10'b0001000010; // 11 * 6 = 66
        rom[359] = 10'b0001001101; // 11 * 7 = 77
        rom[360] = 10'b0001011000; // 11 * 8 = 88
        rom[361] = 10'b0001100011; // 11 * 9 = 99
        rom[362] = 10'b0001101110; // 11 * 10 = 110
        rom[363] = 10'b0001111001; // 11 * 11 = 121
        rom[364] = 10'b0010000100; // 11 * 12 = 132
        rom[365] = 10'b0010001111; // 11 * 13 = 143
        rom[366] = 10'b0010011010; // 11 * 14 = 154
        rom[367] = 10'b0010100101; // 11 * 15 = 165
        rom[368] = 10'b0010110000; // 11 * 16 = 176
        rom[369] = 10'b0010111011; // 11 * 17 = 187
        rom[370] = 10'b0011000110; // 11 * 18 = 198
        rom[371] = 10'b0011010001; // 11 * 19 = 209
        rom[372] = 10'b0011011100; // 11 * 20 = 220
        rom[373] = 10'b0011100111; // 11 * 21 = 231
        rom[374] = 10'b0011110010; // 11 * 22 = 242
        rom[375] = 10'b0011111101; // 11 * 23 = 253
        rom[376] = 10'b0100001000; // 11 * 24 = 264
        rom[377] = 10'b0100010011; // 11 * 25 = 275
        rom[378] = 10'b0100011110; // 11 * 26 = 286
        rom[379] = 10'b0100101001; // 11 * 27 = 297
        rom[380] = 10'b0100110100; // 11 * 28 = 308
        rom[381] = 10'b0100111111; // 11 * 29 = 319
        rom[382] = 10'b0101001010; // 11 * 30 = 330
        rom[383] = 10'b0101010101; // 11 * 31 = 341
        rom[384] = 10'b0000000000; // 12 * 0 = 0
        rom[385] = 10'b0000001100; // 12 * 1 = 12
        rom[386] = 10'b0000011000; // 12 * 2 = 24
        rom[387] = 10'b0000100100; // 12 * 3 = 36
        rom[388] = 10'b0000110000; // 12 * 4 = 48
        rom[389] = 10'b0000111100; // 12 * 5 = 60
        rom[390] = 10'b0001001000; // 12 * 6 = 72
        rom[391] = 10'b0001010100; // 12 * 7 = 84
        rom[392] = 10'b0001100000; // 12 * 8 = 96
        rom[393] = 10'b0001101100; // 12 * 9 = 108
        rom[394] = 10'b0001111000; // 12 * 10 = 120
        rom[395] = 10'b0010000100; // 12 * 11 = 132
        rom[396] = 10'b0010010000; // 12 * 12 = 144
        rom[397] = 10'b0010011100; // 12 * 13 = 156
        rom[398] = 10'b0010101000; // 12 * 14 = 168
        rom[399] = 10'b0010110100; // 12 * 15 = 180
        rom[400] = 10'b0011000000; // 12 * 16 = 192
        rom[401] = 10'b0011001100; // 12 * 17 = 204
        rom[402] = 10'b0011011000; // 12 * 18 = 216
        rom[403] = 10'b0011100100; // 12 * 19 = 228
        rom[404] = 10'b0011110000; // 12 * 20 = 240
        rom[405] = 10'b0011111100; // 12 * 21 = 252
        rom[406] = 10'b0100001000; // 12 * 22 = 264
        rom[407] = 10'b0100010100; // 12 * 23 = 276
        rom[408] = 10'b0100100000; // 12 * 24 = 288
        rom[409] = 10'b0100101100; // 12 * 25 = 300
        rom[410] = 10'b0100111000; // 12 * 26 = 312
        rom[411] = 10'b0101000100; // 12 * 27 = 324
        rom[412] = 10'b0101010000; // 12 * 28 = 336
        rom[413] = 10'b0101011100; // 12 * 29 = 348
        rom[414] = 10'b0101101000; // 12 * 30 = 360
        rom[415] = 10'b0101110100; // 12 * 31 = 372
        rom[416] = 10'b0000000000; // 13 * 0 = 0
        rom[417] = 10'b0000001101; // 13 * 1 = 13
        rom[418] = 10'b0000011010; // 13 * 2 = 26
        rom[419] = 10'b0000100111; // 13 * 3 = 39
        rom[420] = 10'b0000110100; // 13 * 4 = 52
        rom[421] = 10'b0001000001; // 13 * 5 = 65
        rom[422] = 10'b0001001110; // 13 * 6 = 78
        rom[423] = 10'b0001011011; // 13 * 7 = 91
        rom[424] = 10'b0001101000; // 13 * 8 = 104
        rom[425] = 10'b0001110101; // 13 * 9 = 117
        rom[426] = 10'b0010000010; // 13 * 10 = 130
        rom[427] = 10'b0010001111; // 13 * 11 = 143
        rom[428] = 10'b0010011100; // 13 * 12 = 156
        rom[429] = 10'b0010101001; // 13 * 13 = 169
        rom[430] = 10'b0010110110; // 13 * 14 = 182
        rom[431] = 10'b0011000011; // 13 * 15 = 195
        rom[432] = 10'b0011010000; // 13 * 16 = 208
        rom[433] = 10'b0011011101; // 13 * 17 = 221
        rom[434] = 10'b0011101010; // 13 * 18 = 234
        rom[435] = 10'b0011110111; // 13 * 19 = 247
        rom[436] = 10'b0100000100; // 13 * 20 = 260
        rom[437] = 10'b0100010001; // 13 * 21 = 273
        rom[438] = 10'b0100011110; // 13 * 22 = 286
        rom[439] = 10'b0100101011; // 13 * 23 = 299
        rom[440] = 10'b0100111000; // 13 * 24 = 312
        rom[441] = 10'b0101000101; // 13 * 25 = 325
        rom[442] = 10'b0101010010; // 13 * 26 = 338
        rom[443] = 10'b0101011111; // 13 * 27 = 351
        rom[444] = 10'b0101101100; // 13 * 28 = 364
        rom[445] = 10'b0101111001; // 13 * 29 = 377
        rom[446] = 10'b0110000110; // 13 * 30 = 390
        rom[447] = 10'b0110010011; // 13 * 31 = 403
        rom[448] = 10'b0000000000; // 14 * 0 = 0
        rom[449] = 10'b0000001110; // 14 * 1 = 14
        rom[450] = 10'b0000011100; // 14 * 2 = 28
        rom[451] = 10'b0000101010; // 14 * 3 = 42
        rom[452] = 10'b0000111000; // 14 * 4 = 56
        rom[453] = 10'b0001000110; // 14 * 5 = 70
        rom[454] = 10'b0001010100; // 14 * 6 = 84
        rom[455] = 10'b0001100010; // 14 * 7 = 98
        rom[456] = 10'b0001110000; // 14 * 8 = 112
        rom[457] = 10'b0001111110; // 14 * 9 = 126
        rom[458] = 10'b0010001100; // 14 * 10 = 140
        rom[459] = 10'b0010011010; // 14 * 11 = 154
        rom[460] = 10'b0010101000; // 14 * 12 = 168
        rom[461] = 10'b0010110110; // 14 * 13 = 182
        rom[462] = 10'b0011000100; // 14 * 14 = 196
        rom[463] = 10'b0011010010; // 14 * 15 = 210
        rom[464] = 10'b0011100000; // 14 * 16 = 224
        rom[465] = 10'b0011101110; // 14 * 17 = 238
        rom[466] = 10'b0011111100; // 14 * 18 = 252
        rom[467] = 10'b0100001010; // 14 * 19 = 266
        rom[468] = 10'b0100011000; // 14 * 20 = 280
        rom[469] = 10'b0100100110; // 14 * 21 = 294
        rom[470] = 10'b0100110100; // 14 * 22 = 308
        rom[471] = 10'b0101000010; // 14 * 23 = 322
        rom[472] = 10'b0101010000; // 14 * 24 = 336
        rom[473] = 10'b0101011110; // 14 * 25 = 350
        rom[474] = 10'b0101101100; // 14 * 26 = 364
        rom[475] = 10'b0101111010; // 14 * 27 = 378
        rom[476] = 10'b0110001000; // 14 * 28 = 392
        rom[477] = 10'b0110010110; // 14 * 29 = 406
        rom[478] = 10'b0110100100; // 14 * 30 = 420
        rom[479] = 10'b0110110010; // 14 * 31 = 434
        rom[480] = 10'b0000000000; // 15 * 0 = 0
        rom[481] = 10'b0000001111; // 15 * 1 = 15
        rom[482] = 10'b0000011110; // 15 * 2 = 30
        rom[483] = 10'b0000101101; // 15 * 3 = 45
        rom[484] = 10'b0000111100; // 15 * 4 = 60
        rom[485] = 10'b0001001011; // 15 * 5 = 75
        rom[486] = 10'b0001011010; // 15 * 6 = 90
        rom[487] = 10'b0001101001; // 15 * 7 = 105
        rom[488] = 10'b0001111000; // 15 * 8 = 120
        rom[489] = 10'b0010000111; // 15 * 9 = 135
        rom[490] = 10'b0010010110; // 15 * 10 = 150
        rom[491] = 10'b0010100101; // 15 * 11 = 165
        rom[492] = 10'b0010110100; // 15 * 12 = 180
        rom[493] = 10'b0011000011; // 15 * 13 = 195
        rom[494] = 10'b0011010010; // 15 * 14 = 210
        rom[495] = 10'b0011100001; // 15 * 15 = 225
        rom[496] = 10'b0011110000; // 15 * 16 = 240
        rom[497] = 10'b0011111111; // 15 * 17 = 255
        rom[498] = 10'b0100001110; // 15 * 18 = 270
        rom[499] = 10'b0100011101; // 15 * 19 = 285
        rom[500] = 10'b0100101100; // 15 * 20 = 300
        rom[501] = 10'b0100111011; // 15 * 21 = 315
        rom[502] = 10'b0101001010; // 15 * 22 = 330
        rom[503] = 10'b0101011001; // 15 * 23 = 345
        rom[504] = 10'b0101101000; // 15 * 24 = 360
        rom[505] = 10'b0101110111; // 15 * 25 = 375
        rom[506] = 10'b0110000110; // 15 * 26 = 390
        rom[507] = 10'b0110010101; // 15 * 27 = 405
        rom[508] = 10'b0110100100; // 15 * 28 = 420
        rom[509] = 10'b0110110011; // 15 * 29 = 435
        rom[510] = 10'b0111000010; // 15 * 30 = 450
        rom[511] = 10'b0111010001; // 15 * 31 = 465
        rom[512] = 10'b0000000000; // 16 * 0 = 0
        rom[513] = 10'b0000010000; // 16 * 1 = 16
        rom[514] = 10'b0000100000; // 16 * 2 = 32
        rom[515] = 10'b0000110000; // 16 * 3 = 48
        rom[516] = 10'b0001000000; // 16 * 4 = 64
        rom[517] = 10'b0001010000; // 16 * 5 = 80
        rom[518] = 10'b0001100000; // 16 * 6 = 96
        rom[519] = 10'b0001110000; // 16 * 7 = 112
        rom[520] = 10'b0010000000; // 16 * 8 = 128
        rom[521] = 10'b0010010000; // 16 * 9 = 144
        rom[522] = 10'b0010100000; // 16 * 10 = 160
        rom[523] = 10'b0010110000; // 16 * 11 = 176
        rom[524] = 10'b0011000000; // 16 * 12 = 192
        rom[525] = 10'b0011010000; // 16 * 13 = 208
        rom[526] = 10'b0011100000; // 16 * 14 = 224
        rom[527] = 10'b0011110000; // 16 * 15 = 240
        rom[528] = 10'b0100000000; // 16 * 16 = 256
        rom[529] = 10'b0100010000; // 16 * 17 = 272
        rom[530] = 10'b0100100000; // 16 * 18 = 288
        rom[531] = 10'b0100110000; // 16 * 19 = 304
        rom[532] = 10'b0101000000; // 16 * 20 = 320
        rom[533] = 10'b0101010000; // 16 * 21 = 336
        rom[534] = 10'b0101100000; // 16 * 22 = 352
        rom[535] = 10'b0101110000; // 16 * 23 = 368
        rom[536] = 10'b0110000000; // 16 * 24 = 384
        rom[537] = 10'b0110010000; // 16 * 25 = 400
        rom[538] = 10'b0110100000; // 16 * 26 = 416
        rom[539] = 10'b0110110000; // 16 * 27 = 432
        rom[540] = 10'b0111000000; // 16 * 28 = 448
        rom[541] = 10'b0111010000; // 16 * 29 = 464
        rom[542] = 10'b0111100000; // 16 * 30 = 480
        rom[543] = 10'b0111110000; // 16 * 31 = 496
        rom[544] = 10'b0000000000; // 17 * 0 = 0
        rom[545] = 10'b0000010001; // 17 * 1 = 17
        rom[546] = 10'b0000100010; // 17 * 2 = 34
        rom[547] = 10'b0000110011; // 17 * 3 = 51
        rom[548] = 10'b0001000100; // 17 * 4 = 68
        rom[549] = 10'b0001010101; // 17 * 5 = 85
        rom[550] = 10'b0001100110; // 17 * 6 = 102
        rom[551] = 10'b0001110111; // 17 * 7 = 119
        rom[552] = 10'b0010001000; // 17 * 8 = 136
        rom[553] = 10'b0010011001; // 17 * 9 = 153
        rom[554] = 10'b0010101010; // 17 * 10 = 170
        rom[555] = 10'b0010111011; // 17 * 11 = 187
        rom[556] = 10'b0011001100; // 17 * 12 = 204
        rom[557] = 10'b0011011101; // 17 * 13 = 221
        rom[558] = 10'b0011101110; // 17 * 14 = 238
        rom[559] = 10'b0011111111; // 17 * 15 = 255
        rom[560] = 10'b0100010000; // 17 * 16 = 272
        rom[561] = 10'b0100100001; // 17 * 17 = 289
        rom[562] = 10'b0100110010; // 17 * 18 = 306
        rom[563] = 10'b0101000011; // 17 * 19 = 323
        rom[564] = 10'b0101010100; // 17 * 20 = 340
        rom[565] = 10'b0101100101; // 17 * 21 = 357
        rom[566] = 10'b0101110110; // 17 * 22 = 374
        rom[567] = 10'b0110000111; // 17 * 23 = 391
        rom[568] = 10'b0110011000; // 17 * 24 = 408
        rom[569] = 10'b0110101001; // 17 * 25 = 425
        rom[570] = 10'b0110111010; // 17 * 26 = 442
        rom[571] = 10'b0111001011; // 17 * 27 = 459
        rom[572] = 10'b0111011100; // 17 * 28 = 476
        rom[573] = 10'b0111101101; // 17 * 29 = 493
        rom[574] = 10'b0111111110; // 17 * 30 = 510
        rom[575] = 10'b1000001111; // 17 * 31 = 527
        rom[576] = 10'b0000000000; // 18 * 0 = 0
        rom[577] = 10'b0000010010; // 18 * 1 = 18
        rom[578] = 10'b0000100100; // 18 * 2 = 36
        rom[579] = 10'b0000110110; // 18 * 3 = 54
        rom[580] = 10'b0001001000; // 18 * 4 = 72
        rom[581] = 10'b0001011010; // 18 * 5 = 90
        rom[582] = 10'b0001101100; // 18 * 6 = 108
        rom[583] = 10'b0001111110; // 18 * 7 = 126
        rom[584] = 10'b0010010000; // 18 * 8 = 144
        rom[585] = 10'b0010100010; // 18 * 9 = 162
        rom[586] = 10'b0010110100; // 18 * 10 = 180
        rom[587] = 10'b0011000110; // 18 * 11 = 198
        rom[588] = 10'b0011011000; // 18 * 12 = 216
        rom[589] = 10'b0011101010; // 18 * 13 = 234
        rom[590] = 10'b0011111100; // 18 * 14 = 252
        rom[591] = 10'b0100001110; // 18 * 15 = 270
        rom[592] = 10'b0100100000; // 18 * 16 = 288
        rom[593] = 10'b0100110010; // 18 * 17 = 306
        rom[594] = 10'b0101000100; // 18 * 18 = 324
        rom[595] = 10'b0101010110; // 18 * 19 = 342
        rom[596] = 10'b0101101000; // 18 * 20 = 360
        rom[597] = 10'b0101111010; // 18 * 21 = 378
        rom[598] = 10'b0110001100; // 18 * 22 = 396
        rom[599] = 10'b0110011110; // 18 * 23 = 414
        rom[600] = 10'b0110110000; // 18 * 24 = 432
        rom[601] = 10'b0111000010; // 18 * 25 = 450
        rom[602] = 10'b0111010100; // 18 * 26 = 468
        rom[603] = 10'b0111100110; // 18 * 27 = 486
        rom[604] = 10'b0111111000; // 18 * 28 = 504
        rom[605] = 10'b1000001010; // 18 * 29 = 522
        rom[606] = 10'b1000011100; // 18 * 30 = 540
        rom[607] = 10'b1000101110; // 18 * 31 = 558
        rom[608] = 10'b0000000000; // 19 * 0 = 0
        rom[609] = 10'b0000010011; // 19 * 1 = 19
        rom[610] = 10'b0000100110; // 19 * 2 = 38
        rom[611] = 10'b0000111001; // 19 * 3 = 57
        rom[612] = 10'b0001001100; // 19 * 4 = 76
        rom[613] = 10'b0001011111; // 19 * 5 = 95
        rom[614] = 10'b0001110010; // 19 * 6 = 114
        rom[615] = 10'b0010000101; // 19 * 7 = 133
        rom[616] = 10'b0010011000; // 19 * 8 = 152
        rom[617] = 10'b0010101011; // 19 * 9 = 171
        rom[618] = 10'b0010111110; // 19 * 10 = 190
        rom[619] = 10'b0011010001; // 19 * 11 = 209
        rom[620] = 10'b0011100100; // 19 * 12 = 228
        rom[621] = 10'b0011110111; // 19 * 13 = 247
        rom[622] = 10'b0100001010; // 19 * 14 = 266
        rom[623] = 10'b0100011101; // 19 * 15 = 285
        rom[624] = 10'b0100110000; // 19 * 16 = 304
        rom[625] = 10'b0101000011; // 19 * 17 = 323
        rom[626] = 10'b0101010110; // 19 * 18 = 342
        rom[627] = 10'b0101101001; // 19 * 19 = 361
        rom[628] = 10'b0101111100; // 19 * 20 = 380
        rom[629] = 10'b0110001111; // 19 * 21 = 399
        rom[630] = 10'b0110100010; // 19 * 22 = 418
        rom[631] = 10'b0110110101; // 19 * 23 = 437
        rom[632] = 10'b0111001000; // 19 * 24 = 456
        rom[633] = 10'b0111011011; // 19 * 25 = 475
        rom[634] = 10'b0111101110; // 19 * 26 = 494
        rom[635] = 10'b1000000001; // 19 * 27 = 513
        rom[636] = 10'b1000010100; // 19 * 28 = 532
        rom[637] = 10'b1000100111; // 19 * 29 = 551
        rom[638] = 10'b1000111010; // 19 * 30 = 570
        rom[639] = 10'b1001001101; // 19 * 31 = 589
        rom[640] = 10'b0000000000; // 20 * 0 = 0
        rom[641] = 10'b0000010100; // 20 * 1 = 20
        rom[642] = 10'b0000101000; // 20 * 2 = 40
        rom[643] = 10'b0000111100; // 20 * 3 = 60
        rom[644] = 10'b0001010000; // 20 * 4 = 80
        rom[645] = 10'b0001100100; // 20 * 5 = 100
        rom[646] = 10'b0001111000; // 20 * 6 = 120
        rom[647] = 10'b0010001100; // 20 * 7 = 140
        rom[648] = 10'b0010100000; // 20 * 8 = 160
        rom[649] = 10'b0010110100; // 20 * 9 = 180
        rom[650] = 10'b0011001000; // 20 * 10 = 200
        rom[651] = 10'b0011011100; // 20 * 11 = 220
        rom[652] = 10'b0011110000; // 20 * 12 = 240
        rom[653] = 10'b0100000100; // 20 * 13 = 260
        rom[654] = 10'b0100011000; // 20 * 14 = 280
        rom[655] = 10'b0100101100; // 20 * 15 = 300
        rom[656] = 10'b0101000000; // 20 * 16 = 320
        rom[657] = 10'b0101010100; // 20 * 17 = 340
        rom[658] = 10'b0101101000; // 20 * 18 = 360
        rom[659] = 10'b0101111100; // 20 * 19 = 380
        rom[660] = 10'b0110010000; // 20 * 20 = 400
        rom[661] = 10'b0110100100; // 20 * 21 = 420
        rom[662] = 10'b0110111000; // 20 * 22 = 440
        rom[663] = 10'b0111001100; // 20 * 23 = 460
        rom[664] = 10'b0111100000; // 20 * 24 = 480
        rom[665] = 10'b0111110100; // 20 * 25 = 500
        rom[666] = 10'b1000001000; // 20 * 26 = 520
        rom[667] = 10'b1000011100; // 20 * 27 = 540
        rom[668] = 10'b1000110000; // 20 * 28 = 560
        rom[669] = 10'b1001000100; // 20 * 29 = 580
        rom[670] = 10'b1001011000; // 20 * 30 = 600
        rom[671] = 10'b1001101100; // 20 * 31 = 620
        rom[672] = 10'b0000000000; // 21 * 0 = 0
        rom[673] = 10'b0000010101; // 21 * 1 = 21
        rom[674] = 10'b0000101010; // 21 * 2 = 42
        rom[675] = 10'b0000111111; // 21 * 3 = 63
        rom[676] = 10'b0001010100; // 21 * 4 = 84
        rom[677] = 10'b0001101001; // 21 * 5 = 105
        rom[678] = 10'b0001111110; // 21 * 6 = 126
        rom[679] = 10'b0010010011; // 21 * 7 = 147
        rom[680] = 10'b0010101000; // 21 * 8 = 168
        rom[681] = 10'b0010111101; // 21 * 9 = 189
        rom[682] = 10'b0011010010; // 21 * 10 = 210
        rom[683] = 10'b0011100111; // 21 * 11 = 231
        rom[684] = 10'b0011111100; // 21 * 12 = 252
        rom[685] = 10'b0100010001; // 21 * 13 = 273
        rom[686] = 10'b0100100110; // 21 * 14 = 294
        rom[687] = 10'b0100111011; // 21 * 15 = 315
        rom[688] = 10'b0101010000; // 21 * 16 = 336
        rom[689] = 10'b0101100101; // 21 * 17 = 357
        rom[690] = 10'b0101111010; // 21 * 18 = 378
        rom[691] = 10'b0110001111; // 21 * 19 = 399
        rom[692] = 10'b0110100100; // 21 * 20 = 420
        rom[693] = 10'b0110111001; // 21 * 21 = 441
        rom[694] = 10'b0111001110; // 21 * 22 = 462
        rom[695] = 10'b0111100011; // 21 * 23 = 483
        rom[696] = 10'b0111111000; // 21 * 24 = 504
        rom[697] = 10'b1000001101; // 21 * 25 = 525
        rom[698] = 10'b1000100010; // 21 * 26 = 546
        rom[699] = 10'b1000110111; // 21 * 27 = 567
        rom[700] = 10'b1001001100; // 21 * 28 = 588
        rom[701] = 10'b1001100001; // 21 * 29 = 609
        rom[702] = 10'b1001110110; // 21 * 30 = 630
        rom[703] = 10'b1010001011; // 21 * 31 = 651
        rom[704] = 10'b0000000000; // 22 * 0 = 0
        rom[705] = 10'b0000010110; // 22 * 1 = 22
        rom[706] = 10'b0000101100; // 22 * 2 = 44
        rom[707] = 10'b0001000010; // 22 * 3 = 66
        rom[708] = 10'b0001011000; // 22 * 4 = 88
        rom[709] = 10'b0001101110; // 22 * 5 = 110
        rom[710] = 10'b0010000100; // 22 * 6 = 132
        rom[711] = 10'b0010011010; // 22 * 7 = 154
        rom[712] = 10'b0010110000; // 22 * 8 = 176
        rom[713] = 10'b0011000110; // 22 * 9 = 198
        rom[714] = 10'b0011011100; // 22 * 10 = 220
        rom[715] = 10'b0011110010; // 22 * 11 = 242
        rom[716] = 10'b0100001000; // 22 * 12 = 264
        rom[717] = 10'b0100011110; // 22 * 13 = 286
        rom[718] = 10'b0100110100; // 22 * 14 = 308
        rom[719] = 10'b0101001010; // 22 * 15 = 330
        rom[720] = 10'b0101100000; // 22 * 16 = 352
        rom[721] = 10'b0101110110; // 22 * 17 = 374
        rom[722] = 10'b0110001100; // 22 * 18 = 396
        rom[723] = 10'b0110100010; // 22 * 19 = 418
        rom[724] = 10'b0110111000; // 22 * 20 = 440
        rom[725] = 10'b0111001110; // 22 * 21 = 462
        rom[726] = 10'b0111100100; // 22 * 22 = 484
        rom[727] = 10'b0111111010; // 22 * 23 = 506
        rom[728] = 10'b1000010000; // 22 * 24 = 528
        rom[729] = 10'b1000100110; // 22 * 25 = 550
        rom[730] = 10'b1000111100; // 22 * 26 = 572
        rom[731] = 10'b1001010010; // 22 * 27 = 594
        rom[732] = 10'b1001101000; // 22 * 28 = 616
        rom[733] = 10'b1001111110; // 22 * 29 = 638
        rom[734] = 10'b1010010100; // 22 * 30 = 660
        rom[735] = 10'b1010101010; // 22 * 31 = 682
        rom[736] = 10'b0000000000; // 23 * 0 = 0
        rom[737] = 10'b0000010111; // 23 * 1 = 23
        rom[738] = 10'b0000101110; // 23 * 2 = 46
        rom[739] = 10'b0001000101; // 23 * 3 = 69
        rom[740] = 10'b0001011100; // 23 * 4 = 92
        rom[741] = 10'b0001110011; // 23 * 5 = 115
        rom[742] = 10'b0010001010; // 23 * 6 = 138
        rom[743] = 10'b0010100001; // 23 * 7 = 161
        rom[744] = 10'b0010111000; // 23 * 8 = 184
        rom[745] = 10'b0011001111; // 23 * 9 = 207
        rom[746] = 10'b0011100110; // 23 * 10 = 230
        rom[747] = 10'b0011111101; // 23 * 11 = 253
        rom[748] = 10'b0100010100; // 23 * 12 = 276
        rom[749] = 10'b0100101011; // 23 * 13 = 299
        rom[750] = 10'b0101000010; // 23 * 14 = 322
        rom[751] = 10'b0101011001; // 23 * 15 = 345
        rom[752] = 10'b0101110000; // 23 * 16 = 368
        rom[753] = 10'b0110000111; // 23 * 17 = 391
        rom[754] = 10'b0110011110; // 23 * 18 = 414
        rom[755] = 10'b0110110101; // 23 * 19 = 437
        rom[756] = 10'b0111001100; // 23 * 20 = 460
        rom[757] = 10'b0111100011; // 23 * 21 = 483
        rom[758] = 10'b0111111010; // 23 * 22 = 506
        rom[759] = 10'b1000010001; // 23 * 23 = 529
        rom[760] = 10'b1000101000; // 23 * 24 = 552
        rom[761] = 10'b1000111111; // 23 * 25 = 575
        rom[762] = 10'b1001010110; // 23 * 26 = 598
        rom[763] = 10'b1001101101; // 23 * 27 = 621
        rom[764] = 10'b1010000100; // 23 * 28 = 644
        rom[765] = 10'b1010011011; // 23 * 29 = 667
        rom[766] = 10'b1010110010; // 23 * 30 = 690
        rom[767] = 10'b1011001001; // 23 * 31 = 713
        rom[768] = 10'b0000000000; // 24 * 0 = 0
        rom[769] = 10'b0000011000; // 24 * 1 = 24
        rom[770] = 10'b0000110000; // 24 * 2 = 48
        rom[771] = 10'b0001001000; // 24 * 3 = 72
        rom[772] = 10'b0001100000; // 24 * 4 = 96
        rom[773] = 10'b0001111000; // 24 * 5 = 120
        rom[774] = 10'b0010010000; // 24 * 6 = 144
        rom[775] = 10'b0010101000; // 24 * 7 = 168
        rom[776] = 10'b0011000000; // 24 * 8 = 192
        rom[777] = 10'b0011011000; // 24 * 9 = 216
        rom[778] = 10'b0011110000; // 24 * 10 = 240
        rom[779] = 10'b0100001000; // 24 * 11 = 264
        rom[780] = 10'b0100100000; // 24 * 12 = 288
        rom[781] = 10'b0100111000; // 24 * 13 = 312
        rom[782] = 10'b0101010000; // 24 * 14 = 336
        rom[783] = 10'b0101101000; // 24 * 15 = 360
        rom[784] = 10'b0110000000; // 24 * 16 = 384
        rom[785] = 10'b0110011000; // 24 * 17 = 408
        rom[786] = 10'b0110110000; // 24 * 18 = 432
        rom[787] = 10'b0111001000; // 24 * 19 = 456
        rom[788] = 10'b0111100000; // 24 * 20 = 480
        rom[789] = 10'b0111111000; // 24 * 21 = 504
        rom[790] = 10'b1000010000; // 24 * 22 = 528
        rom[791] = 10'b1000101000; // 24 * 23 = 552
        rom[792] = 10'b1001000000; // 24 * 24 = 576
        rom[793] = 10'b1001011000; // 24 * 25 = 600
        rom[794] = 10'b1001110000; // 24 * 26 = 624
        rom[795] = 10'b1010001000; // 24 * 27 = 648
        rom[796] = 10'b1010100000; // 24 * 28 = 672
        rom[797] = 10'b1010111000; // 24 * 29 = 696
        rom[798] = 10'b1011010000; // 24 * 30 = 720
        rom[799] = 10'b1011101000; // 24 * 31 = 744
        rom[800] = 10'b0000000000; // 25 * 0 = 0
        rom[801] = 10'b0000011001; // 25 * 1 = 25
        rom[802] = 10'b0000110010; // 25 * 2 = 50
        rom[803] = 10'b0001001011; // 25 * 3 = 75
        rom[804] = 10'b0001100100; // 25 * 4 = 100
        rom[805] = 10'b0001111101; // 25 * 5 = 125
        rom[806] = 10'b0010010110; // 25 * 6 = 150
        rom[807] = 10'b0010101111; // 25 * 7 = 175
        rom[808] = 10'b0011001000; // 25 * 8 = 200
        rom[809] = 10'b0011100001; // 25 * 9 = 225
        rom[810] = 10'b0011111010; // 25 * 10 = 250
        rom[811] = 10'b0100010011; // 25 * 11 = 275
        rom[812] = 10'b0100101100; // 25 * 12 = 300
        rom[813] = 10'b0101000101; // 25 * 13 = 325
        rom[814] = 10'b0101011110; // 25 * 14 = 350
        rom[815] = 10'b0101110111; // 25 * 15 = 375
        rom[816] = 10'b0110010000; // 25 * 16 = 400
        rom[817] = 10'b0110101001; // 25 * 17 = 425
        rom[818] = 10'b0111000010; // 25 * 18 = 450
        rom[819] = 10'b0111011011; // 25 * 19 = 475
        rom[820] = 10'b0111110100; // 25 * 20 = 500
        rom[821] = 10'b1000001101; // 25 * 21 = 525
        rom[822] = 10'b1000100110; // 25 * 22 = 550
        rom[823] = 10'b1000111111; // 25 * 23 = 575
        rom[824] = 10'b1001011000; // 25 * 24 = 600
        rom[825] = 10'b1001110001; // 25 * 25 = 625
        rom[826] = 10'b1010001010; // 25 * 26 = 650
        rom[827] = 10'b1010100011; // 25 * 27 = 675
        rom[828] = 10'b1010111100; // 25 * 28 = 700
        rom[829] = 10'b1011010101; // 25 * 29 = 725
        rom[830] = 10'b1011101110; // 25 * 30 = 750
        rom[831] = 10'b1100000111; // 25 * 31 = 775
        rom[832] = 10'b0000000000; // 26 * 0 = 0
        rom[833] = 10'b0000011010; // 26 * 1 = 26
        rom[834] = 10'b0000110100; // 26 * 2 = 52
        rom[835] = 10'b0001001110; // 26 * 3 = 78
        rom[836] = 10'b0001101000; // 26 * 4 = 104
        rom[837] = 10'b0010000010; // 26 * 5 = 130
        rom[838] = 10'b0010011100; // 26 * 6 = 156
        rom[839] = 10'b0010110110; // 26 * 7 = 182
        rom[840] = 10'b0011010000; // 26 * 8 = 208
        rom[841] = 10'b0011101010; // 26 * 9 = 234
        rom[842] = 10'b0100000100; // 26 * 10 = 260
        rom[843] = 10'b0100011110; // 26 * 11 = 286
        rom[844] = 10'b0100111000; // 26 * 12 = 312
        rom[845] = 10'b0101010010; // 26 * 13 = 338
        rom[846] = 10'b0101101100; // 26 * 14 = 364
        rom[847] = 10'b0110000110; // 26 * 15 = 390
        rom[848] = 10'b0110100000; // 26 * 16 = 416
        rom[849] = 10'b0110111010; // 26 * 17 = 442
        rom[850] = 10'b0111010100; // 26 * 18 = 468
        rom[851] = 10'b0111101110; // 26 * 19 = 494
        rom[852] = 10'b1000001000; // 26 * 20 = 520
        rom[853] = 10'b1000100010; // 26 * 21 = 546
        rom[854] = 10'b1000111100; // 26 * 22 = 572
        rom[855] = 10'b1001010110; // 26 * 23 = 598
        rom[856] = 10'b1001110000; // 26 * 24 = 624
        rom[857] = 10'b1010001010; // 26 * 25 = 650
        rom[858] = 10'b1010100100; // 26 * 26 = 676
        rom[859] = 10'b1010111110; // 26 * 27 = 702
        rom[860] = 10'b1011011000; // 26 * 28 = 728
        rom[861] = 10'b1011110010; // 26 * 29 = 754
        rom[862] = 10'b1100001100; // 26 * 30 = 780
        rom[863] = 10'b1100100110; // 26 * 31 = 806
        rom[864] = 10'b0000000000; // 27 * 0 = 0
        rom[865] = 10'b0000011011; // 27 * 1 = 27
        rom[866] = 10'b0000110110; // 27 * 2 = 54
        rom[867] = 10'b0001010001; // 27 * 3 = 81
        rom[868] = 10'b0001101100; // 27 * 4 = 108
        rom[869] = 10'b0010000111; // 27 * 5 = 135
        rom[870] = 10'b0010100010; // 27 * 6 = 162
        rom[871] = 10'b0010111101; // 27 * 7 = 189
        rom[872] = 10'b0011011000; // 27 * 8 = 216
        rom[873] = 10'b0011110011; // 27 * 9 = 243
        rom[874] = 10'b0100001110; // 27 * 10 = 270
        rom[875] = 10'b0100101001; // 27 * 11 = 297
        rom[876] = 10'b0101000100; // 27 * 12 = 324
        rom[877] = 10'b0101011111; // 27 * 13 = 351
        rom[878] = 10'b0101111010; // 27 * 14 = 378
        rom[879] = 10'b0110010101; // 27 * 15 = 405
        rom[880] = 10'b0110110000; // 27 * 16 = 432
        rom[881] = 10'b0111001011; // 27 * 17 = 459
        rom[882] = 10'b0111100110; // 27 * 18 = 486
        rom[883] = 10'b1000000001; // 27 * 19 = 513
        rom[884] = 10'b1000011100; // 27 * 20 = 540
        rom[885] = 10'b1000110111; // 27 * 21 = 567
        rom[886] = 10'b1001010010; // 27 * 22 = 594
        rom[887] = 10'b1001101101; // 27 * 23 = 621
        rom[888] = 10'b1010001000; // 27 * 24 = 648
        rom[889] = 10'b1010100011; // 27 * 25 = 675
        rom[890] = 10'b1010111110; // 27 * 26 = 702
        rom[891] = 10'b1011011001; // 27 * 27 = 729
        rom[892] = 10'b1011110100; // 27 * 28 = 756
        rom[893] = 10'b1100001111; // 27 * 29 = 783
        rom[894] = 10'b1100101010; // 27 * 30 = 810
        rom[895] = 10'b1101000101; // 27 * 31 = 837
        rom[896] = 10'b0000000000; // 28 * 0 = 0
        rom[897] = 10'b0000011100; // 28 * 1 = 28
        rom[898] = 10'b0000111000; // 28 * 2 = 56
        rom[899] = 10'b0001010100; // 28 * 3 = 84
        rom[900] = 10'b0001110000; // 28 * 4 = 112
        rom[901] = 10'b0010001100; // 28 * 5 = 140
        rom[902] = 10'b0010101000; // 28 * 6 = 168
        rom[903] = 10'b0011000100; // 28 * 7 = 196
        rom[904] = 10'b0011100000; // 28 * 8 = 224
        rom[905] = 10'b0011111100; // 28 * 9 = 252
        rom[906] = 10'b0100011000; // 28 * 10 = 280
        rom[907] = 10'b0100110100; // 28 * 11 = 308
        rom[908] = 10'b0101010000; // 28 * 12 = 336
        rom[909] = 10'b0101101100; // 28 * 13 = 364
        rom[910] = 10'b0110001000; // 28 * 14 = 392
        rom[911] = 10'b0110100100; // 28 * 15 = 420
        rom[912] = 10'b0111000000; // 28 * 16 = 448
        rom[913] = 10'b0111011100; // 28 * 17 = 476
        rom[914] = 10'b0111111000; // 28 * 18 = 504
        rom[915] = 10'b1000010100; // 28 * 19 = 532
        rom[916] = 10'b1000110000; // 28 * 20 = 560
        rom[917] = 10'b1001001100; // 28 * 21 = 588
        rom[918] = 10'b1001101000; // 28 * 22 = 616
        rom[919] = 10'b1010000100; // 28 * 23 = 644
        rom[920] = 10'b1010100000; // 28 * 24 = 672
        rom[921] = 10'b1010111100; // 28 * 25 = 700
        rom[922] = 10'b1011011000; // 28 * 26 = 728
        rom[923] = 10'b1011110100; // 28 * 27 = 756
        rom[924] = 10'b1100010000; // 28 * 28 = 784
        rom[925] = 10'b1100101100; // 28 * 29 = 812
        rom[926] = 10'b1101001000; // 28 * 30 = 840
        rom[927] = 10'b1101100100; // 28 * 31 = 868
        rom[928] = 10'b0000000000; // 29 * 0 = 0
        rom[929] = 10'b0000011101; // 29 * 1 = 29
        rom[930] = 10'b0000111010; // 29 * 2 = 58
        rom[931] = 10'b0001010111; // 29 * 3 = 87
        rom[932] = 10'b0001110100; // 29 * 4 = 116
        rom[933] = 10'b0010010001; // 29 * 5 = 145
        rom[934] = 10'b0010101110; // 29 * 6 = 174
        rom[935] = 10'b0011001011; // 29 * 7 = 203
        rom[936] = 10'b0011101000; // 29 * 8 = 232
        rom[937] = 10'b0100000101; // 29 * 9 = 261
        rom[938] = 10'b0100100010; // 29 * 10 = 290
        rom[939] = 10'b0100111111; // 29 * 11 = 319
        rom[940] = 10'b0101011100; // 29 * 12 = 348
        rom[941] = 10'b0101111001; // 29 * 13 = 377
        rom[942] = 10'b0110010110; // 29 * 14 = 406
        rom[943] = 10'b0110110011; // 29 * 15 = 435
        rom[944] = 10'b0111010000; // 29 * 16 = 464
        rom[945] = 10'b0111101101; // 29 * 17 = 493
        rom[946] = 10'b1000001010; // 29 * 18 = 522
        rom[947] = 10'b1000100111; // 29 * 19 = 551
        rom[948] = 10'b1001000100; // 29 * 20 = 580
        rom[949] = 10'b1001100001; // 29 * 21 = 609
        rom[950] = 10'b1001111110; // 29 * 22 = 638
        rom[951] = 10'b1010011011; // 29 * 23 = 667
        rom[952] = 10'b1010111000; // 29 * 24 = 696
        rom[953] = 10'b1011010101; // 29 * 25 = 725
        rom[954] = 10'b1011110010; // 29 * 26 = 754
        rom[955] = 10'b1100001111; // 29 * 27 = 783
        rom[956] = 10'b1100101100; // 29 * 28 = 812
        rom[957] = 10'b1101001001; // 29 * 29 = 841
        rom[958] = 10'b1101100110; // 29 * 30 = 870
        rom[959] = 10'b1110000011; // 29 * 31 = 899
        rom[960] = 10'b0000000000; // 30 * 0 = 0
        rom[961] = 10'b0000011110; // 30 * 1 = 30
        rom[962] = 10'b0000111100; // 30 * 2 = 60
        rom[963] = 10'b0001011010; // 30 * 3 = 90
        rom[964] = 10'b0001111000; // 30 * 4 = 120
        rom[965] = 10'b0010010110; // 30 * 5 = 150
        rom[966] = 10'b0010110100; // 30 * 6 = 180
        rom[967] = 10'b0011010010; // 30 * 7 = 210
        rom[968] = 10'b0011110000; // 30 * 8 = 240
        rom[969] = 10'b0100001110; // 30 * 9 = 270
        rom[970] = 10'b0100101100; // 30 * 10 = 300
        rom[971] = 10'b0101001010; // 30 * 11 = 330
        rom[972] = 10'b0101101000; // 30 * 12 = 360
        rom[973] = 10'b0110000110; // 30 * 13 = 390
        rom[974] = 10'b0110100100; // 30 * 14 = 420
        rom[975] = 10'b0111000010; // 30 * 15 = 450
        rom[976] = 10'b0111100000; // 30 * 16 = 480
        rom[977] = 10'b0111111110; // 30 * 17 = 510
        rom[978] = 10'b1000011100; // 30 * 18 = 540
        rom[979] = 10'b1000111010; // 30 * 19 = 570
        rom[980] = 10'b1001011000; // 30 * 20 = 600
        rom[981] = 10'b1001110110; // 30 * 21 = 630
        rom[982] = 10'b1010010100; // 30 * 22 = 660
        rom[983] = 10'b1010110010; // 30 * 23 = 690
        rom[984] = 10'b1011010000; // 30 * 24 = 720
        rom[985] = 10'b1011101110; // 30 * 25 = 750
        rom[986] = 10'b1100001100; // 30 * 26 = 780
        rom[987] = 10'b1100101010; // 30 * 27 = 810
        rom[988] = 10'b1101001000; // 30 * 28 = 840
        rom[989] = 10'b1101100110; // 30 * 29 = 870
        rom[990] = 10'b1110000100; // 30 * 30 = 900
        rom[991] = 10'b1110100010; // 30 * 31 = 930
        rom[992] = 10'b0000000000; // 31 * 0 = 0
        rom[993] = 10'b0000011111; // 31 * 1 = 31
        rom[994] = 10'b0000111110; // 31 * 2 = 62
        rom[995] = 10'b0001011101; // 31 * 3 = 93
        rom[996] = 10'b0001111100; // 31 * 4 = 124
        rom[997] = 10'b0010011011; // 31 * 5 = 155
        rom[998] = 10'b0010111010; // 31 * 6 = 186
        rom[999] = 10'b0011011001; // 31 * 7 = 217
        rom[1000] = 10'b0011111000; // 31 * 8 = 248
        rom[1001] = 10'b0100010111; // 31 * 9 = 279
        rom[1002] = 10'b0100110110; // 31 * 10 = 310
        rom[1003] = 10'b0101010101; // 31 * 11 = 341
        rom[1004] = 10'b0101110100; // 31 * 12 = 372
        rom[1005] = 10'b0110010011; // 31 * 13 = 403
        rom[1006] = 10'b0110110010; // 31 * 14 = 434
        rom[1007] = 10'b0111010001; // 31 * 15 = 465
        rom[1008] = 10'b0111110000; // 31 * 16 = 496
        rom[1009] = 10'b1000001111; // 31 * 17 = 527
        rom[1010] = 10'b1000101110; // 31 * 18 = 558
        rom[1011] = 10'b1001001101; // 31 * 19 = 589
        rom[1012] = 10'b1001101100; // 31 * 20 = 620
        rom[1013] = 10'b1010001011; // 31 * 21 = 651
        rom[1014] = 10'b1010101010; // 31 * 22 = 682
        rom[1015] = 10'b1011001001; // 31 * 23 = 713
        rom[1016] = 10'b1011101000; // 31 * 24 = 744
        rom[1017] = 10'b1100000111; // 31 * 25 = 775
        rom[1018] = 10'b1100100110; // 31 * 26 = 806
        rom[1019] = 10'b1101000101; // 31 * 27 = 837
        rom[1020] = 10'b1101100100; // 31 * 28 = 868
        rom[1021] = 10'b1110000011; // 31 * 29 = 899
        rom[1022] = 10'b1110100010; // 31 * 30 = 930
        rom[1023] = 10'b1111000001; // 31 * 31 = 961

    end

    assign res = rom[{n1,n2}];

endmodule
